module matrixgen(input reset, input clock, input[0:0] address1, input[0:0] address2, input real gate_matrix[0:7], real effective_matrix[0:31]);
  
  parameter NUMBER_OF_QUBITS = 1;
  
endmodule
